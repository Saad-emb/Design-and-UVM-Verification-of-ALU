class env extends uvm_env;
`uvm_component_utils(env)

function new(input string inst = "ENV", uvm_component c);
super.new(inst,c);
endfunction

scoreboard s;
agent a;

virtual function void build_phase(uvm_phase phase);
	super.build_phase(phase);
	a = agent::type_id::create("AGENT",this);
	s = scoreboard::type_id::create("SCO",this);
endfunction

virtual function void connect_phase(uvm_phase phase);
	super.connect_phase(phase);
	//inside monitor send port
	a.m.send.connect(s.recv);
endfunction
endclass
